module genAdder(
	input [4:0] value1,
	input [4:0] value2,
	output [4:0] sum
);

assign sum = value1 + value2;


endmodule