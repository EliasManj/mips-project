module sad_rom_test (

input wire [8:0] addr,
output reg [31:0] dataA,
output reg [31:0] dataB
);

  reg [31:0] rom [0:511];

  always @ * begin
    dataA <= rom[addr];
	  dataB <= rom[addr+256];
  end

  initial begin
  rom[0] = 32'hFFFFFFB7;
  rom[1] = 32'hFFFFFF4E;
  rom[2] = 32'h0000008C;
  rom[3] = 32'hFFFFFF14;
  rom[4] = 32'hFFFFFF2E;
  rom[5] = 32'h0000003D;
  rom[6] = 32'hFFFFFFEE;
  rom[7] = 32'h000000FB;
  rom[8] = 32'hFFFFFF6B;
  rom[9] = 32'hFFFFFFFD;
  rom[10] = 32'hFFFFFF4D;
  rom[11] = 32'hFFFFFF53;
  rom[12] = 32'h000000AD;
  rom[13] = 32'h000000B4;
  rom[14] = 32'hFFFFFFFA;
  rom[15] = 32'h0000008C;
  rom[16] = 32'hFFFFFFB9;
  rom[17] = 32'h0000001E;
  rom[18] = 32'hFFFFFFD9;
  rom[19] = 32'hFFFFFF19;
  rom[20] = 32'hFFFFFF16;
  rom[21] = 32'hFFFFFF3D;
  rom[22] = 32'hFFFFFFAE;
  rom[23] = 32'h00000073;
  rom[24] = 32'hFFFFFF1D;
  rom[25] = 32'h00000057;
  rom[26] = 32'h000000F4;
  rom[27] = 32'h00000030;
  rom[28] = 32'hFFFFFFBD;
  rom[29] = 32'h000000C7;
  rom[30] = 32'h000000F2;
  rom[31] = 32'h000000C5;
  rom[32] = 32'hFFFFFF54;
  rom[33] = 32'hFFFFFF53;
  rom[34] = 32'h0000005E;
  rom[35] = 32'h000000FA;
  rom[36] = 32'hFFFFFF34;
  rom[37] = 32'h00000057;
  rom[38] = 32'hFFFFFF37;
  rom[39] = 32'h000000FE;
  rom[40] = 32'hFFFFFF49;
  rom[41] = 32'hFFFFFF07;
  rom[42] = 32'h000000B0;
  rom[43] = 32'h00000056;
  rom[44] = 32'hFFFFFFBE;
  rom[45] = 32'hFFFFFFDB;
  rom[46] = 32'h00000071;
  rom[47] = 32'h000000F9;
  rom[48] = 32'h00000058;
  rom[49] = 32'hFFFFFF1A;
  rom[50] = 32'h000000C4;
  rom[51] = 32'h00000031;
  rom[52] = 32'h00000028;
  rom[53] = 32'hFFFFFFF2;
  rom[54] = 32'h00000028;
  rom[55] = 32'hFFFFFFBC;
  rom[56] = 32'h0000001A;
  rom[57] = 32'h000000D1;
  rom[58] = 32'h0000007A;
  rom[59] = 32'hFFFFFF28;
  rom[60] = 32'h000000C9;
  rom[61] = 32'h000000BE;
  rom[62] = 32'hFFFFFF4D;
  rom[63] = 32'hFFFFFFC3;
  rom[64] = 32'h000000DF;
  rom[65] = 32'h000000D6;
  rom[66] = 32'hFFFFFF28;
  rom[67] = 32'h0000007E;
  rom[68] = 32'hFFFFFF17;
  rom[69] = 32'h00000004;
  rom[70] = 32'hFFFFFF2F;
  rom[71] = 32'hFFFFFF72;
  rom[72] = 32'hFFFFFF1C;
  rom[73] = 32'h000000DA;
  rom[74] = 32'h000000D7;
  rom[75] = 32'hFFFFFF4F;
  rom[76] = 32'hFFFFFFEA;
  rom[77] = 32'h00000003;
  rom[78] = 32'hFFFFFF1D;
  rom[79] = 32'h00000003;
  rom[80] = 32'h0000001E;
  rom[81] = 32'hFFFFFF07;
  rom[82] = 32'hFFFFFF7E;
  rom[83] = 32'hFFFFFFAC;
  rom[84] = 32'h00000079;
  rom[85] = 32'h00000004;
  rom[86] = 32'h000000CB;
  rom[87] = 32'h00000097;
  rom[88] = 32'hFFFFFF1D;
  rom[89] = 32'h00000074;
  rom[90] = 32'h0000008D;
  rom[91] = 32'h00000031;
  rom[92] = 32'h0000002A;
  rom[93] = 32'hFFFFFF2D;
  rom[94] = 32'hFFFFFF16;
  rom[95] = 32'hFFFFFFC5;
  rom[96] = 32'hFFFFFFAC;
  rom[97] = 32'h000000F4;
  rom[98] = 32'hFFFFFFFA;
  rom[99] = 32'h000000FB;
  rom[100] = 32'h000000AD;
  rom[101] = 32'h000000FD;
  rom[102] = 32'hFFFFFF50;
  rom[103] = 32'hFFFFFFA7;
  rom[104] = 32'hFFFFFFD8;
  rom[105] = 32'hFFFFFF59;
  rom[106] = 32'hFFFFFF87;
  rom[107] = 32'h00000045;
  rom[108] = 32'hFFFFFF4B;
  rom[109] = 32'h00000079;
  rom[110] = 32'h000000A4;
  rom[111] = 32'hFFFFFF2D;
  rom[112] = 32'hFFFFFF0F;
  rom[113] = 32'hFFFFFF7C;
  rom[114] = 32'h000000AC;
  rom[115] = 32'h0000005A;
  rom[116] = 32'hFFFFFF76;
  rom[117] = 32'h000000FE;
  rom[118] = 32'hFFFFFF92;
  rom[119] = 32'hFFFFFFA4;
  rom[120] = 32'h00000076;
  rom[121] = 32'h00000065;
  rom[122] = 32'hFFFFFF35;
  rom[123] = 32'h00000040;
  rom[124] = 32'hFFFFFF26;
  rom[125] = 32'hFFFFFFF9;
  rom[126] = 32'hFFFFFFD8;
  rom[127] = 32'hFFFFFFD2;
  rom[128] = 32'hFFFFFF8A;
  rom[129] = 32'hFFFFFF61;
  rom[130] = 32'hFFFFFFE6;
  rom[131] = 32'hFFFFFF0C;
  rom[132] = 32'h000000B9;
  rom[133] = 32'h00000032;
  rom[134] = 32'hFFFFFF15;
  rom[135] = 32'hFFFFFFAA;
  rom[136] = 32'hFFFFFFF7;
  rom[137] = 32'hFFFFFF4F;
  rom[138] = 32'h000000B7;
  rom[139] = 32'h00000021;
  rom[140] = 32'hFFFFFFD3;
  rom[141] = 32'h0000005D;
  rom[142] = 32'hFFFFFF40;
  rom[143] = 32'h000000BC;
  rom[144] = 32'h0000001E;
  rom[145] = 32'h0000004D;
  rom[146] = 32'h00000054;
  rom[147] = 32'h00000014;
  rom[148] = 32'h000000C3;
  rom[149] = 32'h0000008F;
  rom[150] = 32'hFFFFFF32;
  rom[151] = 32'h00000087;
  rom[152] = 32'h00000077;
  rom[153] = 32'hFFFFFFAE;
  rom[154] = 32'hFFFFFFC1;
  rom[155] = 32'h00000099;
  rom[156] = 32'h0000005A;
  rom[157] = 32'hFFFFFF54;
  rom[158] = 32'h0000001A;
  rom[159] = 32'h0000007F;
  rom[160] = 32'hFFFFFF3D;
  rom[161] = 32'h00000040;
  rom[162] = 32'h000000A0;
  rom[163] = 32'h000000C1;
  rom[164] = 32'h00000047;
  rom[165] = 32'h00000034;
  rom[166] = 32'hFFFFFF2A;
  rom[167] = 32'h00000044;
  rom[168] = 32'h000000F8;
  rom[169] = 32'hFFFFFFC9;
  rom[170] = 32'h00000072;
  rom[171] = 32'hFFFFFFF7;
  rom[172] = 32'h00000045;
  rom[173] = 32'hFFFFFFAF;
  rom[174] = 32'hFFFFFF4E;
  rom[175] = 32'hFFFFFF50;
  rom[176] = 32'hFFFFFF16;
  rom[177] = 32'hFFFFFF2D;
  rom[178] = 32'h0000007F;
  rom[179] = 32'hFFFFFFAC;
  rom[180] = 32'h000000D1;
  rom[181] = 32'h00000013;
  rom[182] = 32'hFFFFFF1B;
  rom[183] = 32'hFFFFFF46;
  rom[184] = 32'hFFFFFFE8;
  rom[185] = 32'h00000064;
  rom[186] = 32'hFFFFFFE2;
  rom[187] = 32'hFFFFFF2C;
  rom[188] = 32'hFFFFFF23;
  rom[189] = 32'hFFFFFF08;
  rom[190] = 32'hFFFFFFA6;
  rom[191] = 32'h000000A2;
  rom[192] = 32'h000000BF;
  rom[193] = 32'h000000E9;
  rom[194] = 32'h000000FB;
  rom[195] = 32'hFFFFFF10;
  rom[196] = 32'hFFFFFF6C;
  rom[197] = 32'hFFFFFF74;
  rom[198] = 32'h00000049;
  rom[199] = 32'hFFFFFFC2;
  rom[200] = 32'hFFFFFF57;
  rom[201] = 32'hFFFFFFA6;
  rom[202] = 32'h00000008;
  rom[203] = 32'hFFFFFF30;
  rom[204] = 32'h000000CB;
  rom[205] = 32'h000000F3;
  rom[206] = 32'h00000033;
  rom[207] = 32'h00000063;
  rom[208] = 32'h00000004;
  rom[209] = 32'h00000060;
  rom[210] = 32'hFFFFFF0D;
  rom[211] = 32'h0000008D;
  rom[212] = 32'hFFFFFF42;
  rom[213] = 32'h000000D8;
  rom[214] = 32'hFFFFFFCC;
  rom[215] = 32'hFFFFFFC5;
  rom[216] = 32'hFFFFFFE2;
  rom[217] = 32'hFFFFFFEA;
  rom[218] = 32'h000000F7;
  rom[219] = 32'h0000008A;
  rom[220] = 32'hFFFFFF9E;
  rom[221] = 32'hFFFFFF9A;
  rom[222] = 32'h000000BF;
  rom[223] = 32'h000000D8;
  rom[224] = 32'hFFFFFF93;
  rom[225] = 32'h000000C9;
  rom[226] = 32'hFFFFFFA9;
  rom[227] = 32'h00000054;
  rom[228] = 32'h000000FD;
  rom[229] = 32'h000000C6;
  rom[230] = 32'hFFFFFF33;
  rom[231] = 32'hFFFFFFFF;
  rom[232] = 32'h000000EF;
  rom[233] = 32'h00000017;
  rom[234] = 32'hFFFFFF22;
  rom[235] = 32'hFFFFFFE4;
  rom[236] = 32'hFFFFFFE2;
  rom[237] = 32'h000000FE;
  rom[238] = 32'hFFFFFF4D;
  rom[239] = 32'hFFFFFFD0;
  rom[240] = 32'hFFFFFF6B;
  rom[241] = 32'hFFFFFF8A;
  rom[242] = 32'hFFFFFFCC;
  rom[243] = 32'h00000010;
  rom[244] = 32'hFFFFFF6D;
  rom[245] = 32'hFFFFFFBE;
  rom[246] = 32'h00000029;
  rom[247] = 32'hFFFFFF47;
  rom[248] = 32'hFFFFFFCA;
  rom[249] = 32'hFFFFFF42;
  rom[250] = 32'hFFFFFF8C;
  rom[251] = 32'hFFFFFF25;
  rom[252] = 32'h00000020;
  rom[253] = 32'hFFFFFF5A;
  rom[254] = 32'h00000073;
  rom[255] = 32'hFFFFFF16;
  rom[256] = 32'h000000D5;
  rom[257] = 32'hFFFFFFF0;
  rom[258] = 32'hFFFFFF3F;
  rom[259] = 32'h000000A0;
  rom[260] = 32'hFFFFFF7A;
  rom[261] = 32'h000000BA;
  rom[262] = 32'h0000006E;
  rom[263] = 32'hFFFFFF17;
  rom[264] = 32'hFFFFFF4D;
  rom[265] = 32'hFFFFFFE3;
  rom[266] = 32'hFFFFFF6C;
  rom[267] = 32'hFFFFFF66;
  rom[268] = 32'h000000E5;
  rom[269] = 32'h0000006E;
  rom[270] = 32'h000000F4;
  rom[271] = 32'hFFFFFFBE;
  rom[272] = 32'h000000B9;
  rom[273] = 32'hFFFFFF8D;
  rom[274] = 32'hFFFFFF49;
  rom[275] = 32'h00000043;
  rom[276] = 32'h000000ED;
  rom[277] = 32'h0000005B;
  rom[278] = 32'h0000008F;
  rom[279] = 32'hFFFFFFBC;
  rom[280] = 32'h00000048;
  rom[281] = 32'hFFFFFF0E;
  rom[282] = 32'h00000033;
  rom[283] = 32'hFFFFFFD3;
  rom[284] = 32'hFFFFFF0E;
  rom[285] = 32'hFFFFFF3C;
  rom[286] = 32'hFFFFFF30;
  rom[287] = 32'hFFFFFFC6;
  rom[288] = 32'hFFFFFF84;
  rom[289] = 32'h00000014;
  rom[290] = 32'hFFFFFF4A;
  rom[291] = 32'hFFFFFFE0;
  rom[292] = 32'h00000039;
  rom[293] = 32'hFFFFFF7F;
  rom[294] = 32'h00000000;
  rom[295] = 32'h00000036;
  rom[296] = 32'hFFFFFF98;
  rom[297] = 32'hFFFFFFDC;
  rom[298] = 32'h000000CE;
  rom[299] = 32'h0000002D;
  rom[300] = 32'hFFFFFFCB;
  rom[301] = 32'hFFFFFFAC;
  rom[302] = 32'hFFFFFF4A;
  rom[303] = 32'h0000000C;
  rom[304] = 32'h000000FB;
  rom[305] = 32'h00000055;
  rom[306] = 32'hFFFFFF07;
  rom[307] = 32'h0000006C;
  rom[308] = 32'h0000006A;
  rom[309] = 32'hFFFFFF2A;
  rom[310] = 32'h00000012;
  rom[311] = 32'h00000060;
  rom[312] = 32'h0000000A;
  rom[313] = 32'hFFFFFFD3;
  rom[314] = 32'hFFFFFF16;
  rom[315] = 32'h0000008D;
  rom[316] = 32'hFFFFFFDA;
  rom[317] = 32'hFFFFFFAF;
  rom[318] = 32'hFFFFFF35;
  rom[319] = 32'hFFFFFFBC;
  rom[320] = 32'h00000087;
  rom[321] = 32'h0000007D;
  rom[322] = 32'h0000003A;
  rom[323] = 32'hFFFFFFAA;
  rom[324] = 32'h00000023;
  rom[325] = 32'hFFFFFFA8;
  rom[326] = 32'hFFFFFF19;
  rom[327] = 32'h00000081;
  rom[328] = 32'h00000065;
  rom[329] = 32'hFFFFFFDA;
  rom[330] = 32'hFFFFFFAB;
  rom[331] = 32'hFFFFFFF8;
  rom[332] = 32'h00000093;
  rom[333] = 32'hFFFFFFBB;
  rom[334] = 32'hFFFFFFB7;
  rom[335] = 32'h000000A5;
  rom[336] = 32'h00000000;
  rom[337] = 32'hFFFFFF0E;
  rom[338] = 32'h00000016;
  rom[339] = 32'hFFFFFF1F;
  rom[340] = 32'hFFFFFF26;
  rom[341] = 32'hFFFFFF59;
  rom[342] = 32'h00000075;
  rom[343] = 32'h00000063;
  rom[344] = 32'hFFFFFF66;
  rom[345] = 32'hFFFFFF93;
  rom[346] = 32'h000000BD;
  rom[347] = 32'hFFFFFF67;
  rom[348] = 32'h000000B4;
  rom[349] = 32'h00000071;
  rom[350] = 32'hFFFFFF75;
  rom[351] = 32'h00000067;
  rom[352] = 32'h0000008E;
  rom[353] = 32'hFFFFFF2F;
  rom[354] = 32'h0000003F;
  rom[355] = 32'h00000050;
  rom[356] = 32'h00000026;
  rom[357] = 32'h00000023;
  rom[358] = 32'hFFFFFF0B;
  rom[359] = 32'h000000D2;
  rom[360] = 32'h00000083;
  rom[361] = 32'h000000C0;
  rom[362] = 32'h00000079;
  rom[363] = 32'h00000060;
  rom[364] = 32'hFFFFFF4F;
  rom[365] = 32'h0000003B;
  rom[366] = 32'h00000036;
  rom[367] = 32'h000000FE;
  rom[368] = 32'hFFFFFFB0;
  rom[369] = 32'hFFFFFF95;
  rom[370] = 32'hFFFFFF0B;
  rom[371] = 32'h000000A8;
  rom[372] = 32'hFFFFFF7D;
  rom[373] = 32'hFFFFFF97;
  rom[374] = 32'hFFFFFF33;
  rom[375] = 32'h0000009A;
  rom[376] = 32'h000000BA;
  rom[377] = 32'h0000003F;
  rom[378] = 32'h00000080;
  rom[379] = 32'h00000069;
  rom[380] = 32'hFFFFFF35;
  rom[381] = 32'h0000002A;
  rom[382] = 32'h00000093;
  rom[383] = 32'hFFFFFF54;
  rom[384] = 32'h00000023;
  rom[385] = 32'h00000088;
  rom[386] = 32'h00000048;
  rom[387] = 32'hFFFFFF0E;
  rom[388] = 32'hFFFFFFFE;
  rom[389] = 32'hFFFFFF71;
  rom[390] = 32'h0000004E;
  rom[391] = 32'hFFFFFF75;
  rom[392] = 32'hFFFFFFBE;
  rom[393] = 32'h000000CC;
  rom[394] = 32'hFFFFFF2C;
  rom[395] = 32'h00000083;
  rom[396] = 32'h0000005B;
  rom[397] = 32'h0000004C;
  rom[398] = 32'hFFFFFF73;
  rom[399] = 32'hFFFFFF45;
  rom[400] = 32'hFFFFFF07;
  rom[401] = 32'h0000000B;
  rom[402] = 32'h000000A6;
  rom[403] = 32'h0000006C;
  rom[404] = 32'h0000007E;
  rom[405] = 32'hFFFFFFD5;
  rom[406] = 32'h0000004A;
  rom[407] = 32'hFFFFFF92;
  rom[408] = 32'hFFFFFF40;
  rom[409] = 32'h0000003C;
  rom[410] = 32'h00000046;
  rom[411] = 32'hFFFFFF49;
  rom[412] = 32'h00000095;
  rom[413] = 32'h000000AF;
  rom[414] = 32'hFFFFFFE1;
  rom[415] = 32'hFFFFFF0A;
  rom[416] = 32'hFFFFFFB3;
  rom[417] = 32'h0000006E;
  rom[418] = 32'h000000C0;
  rom[419] = 32'h00000084;
  rom[420] = 32'h00000014;
  rom[421] = 32'hFFFFFF48;
  rom[422] = 32'h000000C1;
  rom[423] = 32'hFFFFFF0D;
  rom[424] = 32'h000000A7;
  rom[425] = 32'h00000015;
  rom[426] = 32'hFFFFFFD2;
  rom[427] = 32'hFFFFFF5E;
  rom[428] = 32'h000000DD;
  rom[429] = 32'hFFFFFFA2;
  rom[430] = 32'hFFFFFF7C;
  rom[431] = 32'h00000080;
  rom[432] = 32'h00000060;
  rom[433] = 32'h00000090;
  rom[434] = 32'hFFFFFFB4;
  rom[435] = 32'h000000E0;
  rom[436] = 32'hFFFFFFFC;
  rom[437] = 32'h00000073;
  rom[438] = 32'hFFFFFF96;
  rom[439] = 32'hFFFFFF52;
  rom[440] = 32'h000000CA;
  rom[441] = 32'h000000FA;
  rom[442] = 32'hFFFFFF61;
  rom[443] = 32'h000000E7;
  rom[444] = 32'h00000078;
  rom[445] = 32'hFFFFFFEE;
  rom[446] = 32'hFFFFFFD4;
  rom[447] = 32'h0000000E;
  rom[448] = 32'hFFFFFF94;
  rom[449] = 32'h00000034;
  rom[450] = 32'h000000C0;
  rom[451] = 32'h00000087;
  rom[452] = 32'h0000008E;
  rom[453] = 32'hFFFFFF1A;
  rom[454] = 32'h00000064;
  rom[455] = 32'hFFFFFFDA;
  rom[456] = 32'h00000045;
  rom[457] = 32'h00000039;
  rom[458] = 32'hFFFFFFE3;
  rom[459] = 32'h0000005C;
  rom[460] = 32'hFFFFFF9D;
  rom[461] = 32'hFFFFFFFE;
  rom[462] = 32'hFFFFFF8F;
  rom[463] = 32'hFFFFFF62;
  rom[464] = 32'h00000039;
  rom[465] = 32'hFFFFFF32;
  rom[466] = 32'h00000032;
  rom[467] = 32'h000000E5;
  rom[468] = 32'h0000008E;
  rom[469] = 32'hFFFFFF7D;
  rom[470] = 32'hFFFFFF5F;
  rom[471] = 32'h00000071;
  rom[472] = 32'h00000028;
  rom[473] = 32'h00000098;
  rom[474] = 32'hFFFFFF4B;
  rom[475] = 32'hFFFFFF06;
  rom[476] = 32'h00000069;
  rom[477] = 32'h00000079;
  rom[478] = 32'h000000A2;
  rom[479] = 32'h00000037;
  rom[480] = 32'h000000C5;
  rom[481] = 32'h0000009F;
  rom[482] = 32'hFFFFFF57;
  rom[483] = 32'hFFFFFFF0;
  rom[484] = 32'h000000BA;
  rom[485] = 32'h000000FD;
  rom[486] = 32'h000000BA;
  rom[487] = 32'h00000075;
  rom[488] = 32'h0000003B;
  rom[489] = 32'hFFFFFFD8;
  rom[490] = 32'h000000E3;
  rom[491] = 32'hFFFFFF6E;
  rom[492] = 32'h0000000B;
  rom[493] = 32'hFFFFFF9C;
  rom[494] = 32'h00000019;
  rom[495] = 32'h000000BB;
  rom[496] = 32'hFFFFFF92;
  rom[497] = 32'hFFFFFF39;
  rom[498] = 32'h000000FE;
  rom[499] = 32'h0000004D;
  rom[500] = 32'h00000070;
  rom[501] = 32'h0000008F;
  rom[502] = 32'hFFFFFF9A;
  rom[503] = 32'hFFFFFF4D;
  rom[504] = 32'hFFFFFFE9;
  rom[505] = 32'hFFFFFF7D;
  rom[506] = 32'h00000000;
  rom[507] = 32'h00000071;
  rom[508] = 32'h000000D6;
  rom[509] = 32'hFFFFFF05;
  rom[510] = 32'hFFFFFF58;
  rom[511] = 32'hFFFFFF84;

   end
endmodule
