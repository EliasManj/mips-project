module genram2 #(             //-- Parametros
         parameter AW = 9,   //-- Bits de las direcciones (Adress width)
         parameter DW = 32	)   //-- Bits de los datos (Data witdh)

       (        //-- Puertos
         input clk,                      //-- Se�al de reloj global
         input wire [AW-1: 0] addr,      //-- Direcciones
         input wire rw,                  //-- Modo lectura (1) o escritura (0)
         input wire [DW-1: 0] data_in,   //-- Dato de entrada
         output reg [DW-1: 0] data_out); //-- Dato a escribir

//-- Parametro: Nombre del fichero con el contenido de la RAM



//-- Calcular el numero de posiciones totales de memoria
localparam NPOS = 2 ** AW;

  //-- Memoria
  reg [DW-1: 0] ram [0: NPOS-1];

initial begin
ram[0] = 32'hFFFFFFB7;
ram[1] = 32'hFFFFFF4E;
ram[2] = 32'h0000008C;
ram[3] = 32'hFFFFFF14;
ram[4] = 32'hFFFFFF2E;
ram[5] = 32'h0000003D;
ram[6] = 32'hFFFFFFEE;
ram[7] = 32'h000000FB;
ram[8] = 32'hFFFFFF6B;
ram[9] = 32'hFFFFFFFD;
ram[10] = 32'hFFFFFF4D;
ram[11] = 32'hFFFFFF53;
ram[12] = 32'h000000AD;
ram[13] = 32'h000000B4;
ram[14] = 32'hFFFFFFFA;
ram[15] = 32'h0000008C;
ram[16] = 32'hFFFFFFB9;
ram[17] = 32'h0000001E;
ram[18] = 32'hFFFFFFD9;
ram[19] = 32'hFFFFFF19;
ram[20] = 32'hFFFFFF16;
ram[21] = 32'hFFFFFF3D;
ram[22] = 32'hFFFFFFAE;
ram[23] = 32'h00000073;
ram[24] = 32'hFFFFFF1D;
ram[25] = 32'h00000057;
ram[26] = 32'h000000F4;
ram[27] = 32'h00000030;
ram[28] = 32'hFFFFFFBD;
ram[29] = 32'h000000C7;
ram[30] = 32'h000000F2;
ram[31] = 32'h000000C5;
ram[32] = 32'hFFFFFF54;
ram[33] = 32'hFFFFFF53;
ram[34] = 32'h0000005E;
ram[35] = 32'h000000FA;
ram[36] = 32'hFFFFFF34;
ram[37] = 32'h00000057;
ram[38] = 32'hFFFFFF37;
ram[39] = 32'h000000FE;
ram[40] = 32'hFFFFFF49;
ram[41] = 32'hFFFFFF07;
ram[42] = 32'h000000B0;
ram[43] = 32'h00000056;
ram[44] = 32'hFFFFFFBE;
ram[45] = 32'hFFFFFFDB;
ram[46] = 32'h00000071;
ram[47] = 32'h000000F9;
ram[48] = 32'h00000058;
ram[49] = 32'hFFFFFF1A;
ram[50] = 32'h000000C4;
ram[51] = 32'h00000031;
ram[52] = 32'h00000028;
ram[53] = 32'hFFFFFFF2;
ram[54] = 32'h00000028;
ram[55] = 32'hFFFFFFBC;
ram[56] = 32'h0000001A;
ram[57] = 32'h000000D1;
ram[58] = 32'h0000007A;
ram[59] = 32'hFFFFFF28;
ram[60] = 32'h000000C9;
ram[61] = 32'h000000BE;
ram[62] = 32'hFFFFFF4D;
ram[63] = 32'hFFFFFFC3;
ram[64] = 32'h000000DF;
ram[65] = 32'h000000D6;
ram[66] = 32'hFFFFFF28;
ram[67] = 32'h0000007E;
ram[68] = 32'hFFFFFF17;
ram[69] = 32'h00000004;
ram[70] = 32'hFFFFFF2F;
ram[71] = 32'hFFFFFF72;
ram[72] = 32'hFFFFFF1C;
ram[73] = 32'h000000DA;
ram[74] = 32'h000000D7;
ram[75] = 32'hFFFFFF4F;
ram[76] = 32'hFFFFFFEA;
ram[77] = 32'h00000003;
ram[78] = 32'hFFFFFF1D;
ram[79] = 32'h00000003;
ram[80] = 32'h0000001E;
ram[81] = 32'hFFFFFF07;
ram[82] = 32'hFFFFFF7E;
ram[83] = 32'hFFFFFFAC;
ram[84] = 32'h00000079;
ram[85] = 32'h00000004;
ram[86] = 32'h000000CB;
ram[87] = 32'h00000097;
ram[88] = 32'hFFFFFF1D;
ram[89] = 32'h00000074;
ram[90] = 32'h0000008D;
ram[91] = 32'h00000031;
ram[92] = 32'h0000002A;
ram[93] = 32'hFFFFFF2D;
ram[94] = 32'hFFFFFF16;
ram[95] = 32'hFFFFFFC5;
ram[96] = 32'hFFFFFFAC;
ram[97] = 32'h000000F4;
ram[98] = 32'hFFFFFFFA;
ram[99] = 32'h000000FB;
ram[100] = 32'h000000AD;
ram[101] = 32'h000000FD;
ram[102] = 32'hFFFFFF50;
ram[103] = 32'hFFFFFFA7;
ram[104] = 32'hFFFFFFD8;
ram[105] = 32'hFFFFFF59;
ram[106] = 32'hFFFFFF87;
ram[107] = 32'h00000045;
ram[108] = 32'hFFFFFF4B;
ram[109] = 32'h00000079;
ram[110] = 32'h000000A4;
ram[111] = 32'hFFFFFF2D;
ram[112] = 32'hFFFFFF0F;
ram[113] = 32'hFFFFFF7C;
ram[114] = 32'h000000AC;
ram[115] = 32'h0000005A;
ram[116] = 32'hFFFFFF76;
ram[117] = 32'h000000FE;
ram[118] = 32'hFFFFFF92;
ram[119] = 32'hFFFFFFA4;
ram[120] = 32'h00000076;
ram[121] = 32'h00000065;
ram[122] = 32'hFFFFFF35;
ram[123] = 32'h00000040;
ram[124] = 32'hFFFFFF26;
ram[125] = 32'hFFFFFFF9;
ram[126] = 32'hFFFFFFD8;
ram[127] = 32'hFFFFFFD2;
ram[128] = 32'hFFFFFF8A;
ram[129] = 32'hFFFFFF61;
ram[130] = 32'hFFFFFFE6;
ram[131] = 32'hFFFFFF0C;
ram[132] = 32'h000000B9;
ram[133] = 32'h00000032;
ram[134] = 32'hFFFFFF15;
ram[135] = 32'hFFFFFFAA;
ram[136] = 32'hFFFFFFF7;
ram[137] = 32'hFFFFFF4F;
ram[138] = 32'h000000B7;
ram[139] = 32'h00000021;
ram[140] = 32'hFFFFFFD3;
ram[141] = 32'h0000005D;
ram[142] = 32'hFFFFFF40;
ram[143] = 32'h000000BC;
ram[144] = 32'h0000001E;
ram[145] = 32'h0000004D;
ram[146] = 32'h00000054;
ram[147] = 32'h00000014;
ram[148] = 32'h000000C3;
ram[149] = 32'h0000008F;
ram[150] = 32'hFFFFFF32;
ram[151] = 32'h00000087;
ram[152] = 32'h00000077;
ram[153] = 32'hFFFFFFAE;
ram[154] = 32'hFFFFFFC1;
ram[155] = 32'h00000099;
ram[156] = 32'h0000005A;
ram[157] = 32'hFFFFFF54;
ram[158] = 32'h0000001A;
ram[159] = 32'h0000007F;
ram[160] = 32'hFFFFFF3D;
ram[161] = 32'h00000040;
ram[162] = 32'h000000A0;
ram[163] = 32'h000000C1;
ram[164] = 32'h00000047;
ram[165] = 32'h00000034;
ram[166] = 32'hFFFFFF2A;
ram[167] = 32'h00000044;
ram[168] = 32'h000000F8;
ram[169] = 32'hFFFFFFC9;
ram[170] = 32'h00000072;
ram[171] = 32'hFFFFFFF7;
ram[172] = 32'h00000045;
ram[173] = 32'hFFFFFFAF;
ram[174] = 32'hFFFFFF4E;
ram[175] = 32'hFFFFFF50;
ram[176] = 32'hFFFFFF16;
ram[177] = 32'hFFFFFF2D;
ram[178] = 32'h0000007F;
ram[179] = 32'hFFFFFFAC;
ram[180] = 32'h000000D1;
ram[181] = 32'h00000013;
ram[182] = 32'hFFFFFF1B;
ram[183] = 32'hFFFFFF46;
ram[184] = 32'hFFFFFFE8;
ram[185] = 32'h00000064;
ram[186] = 32'hFFFFFFE2;
ram[187] = 32'hFFFFFF2C;
ram[188] = 32'hFFFFFF23;
ram[189] = 32'hFFFFFF08;
ram[190] = 32'hFFFFFFA6;
ram[191] = 32'h000000A2;
ram[192] = 32'h000000BF;
ram[193] = 32'h000000E9;
ram[194] = 32'h000000FB;
ram[195] = 32'hFFFFFF10;
ram[196] = 32'hFFFFFF6C;
ram[197] = 32'hFFFFFF74;
ram[198] = 32'h00000049;
ram[199] = 32'hFFFFFFC2;
ram[200] = 32'hFFFFFF57;
ram[201] = 32'hFFFFFFA6;
ram[202] = 32'h00000008;
ram[203] = 32'hFFFFFF30;
ram[204] = 32'h000000CB;
ram[205] = 32'h000000F3;
ram[206] = 32'h00000033;
ram[207] = 32'h00000063;
ram[208] = 32'h00000004;
ram[209] = 32'h00000060;
ram[210] = 32'hFFFFFF0D;
ram[211] = 32'h0000008D;
ram[212] = 32'hFFFFFF42;
ram[213] = 32'h000000D8;
ram[214] = 32'hFFFFFFCC;
ram[215] = 32'hFFFFFFC5;
ram[216] = 32'hFFFFFFE2;
ram[217] = 32'hFFFFFFEA;
ram[218] = 32'h000000F7;
ram[219] = 32'h0000008A;
ram[220] = 32'hFFFFFF9E;
ram[221] = 32'hFFFFFF9A;
ram[222] = 32'h000000BF;
ram[223] = 32'h000000D8;
ram[224] = 32'hFFFFFF93;
ram[225] = 32'h000000C9;
ram[226] = 32'hFFFFFFA9;
ram[227] = 32'h00000054;
ram[228] = 32'h000000FD;
ram[229] = 32'h000000C6;
ram[230] = 32'hFFFFFF33;
ram[231] = 32'hFFFFFFFF;
ram[232] = 32'h000000EF;
ram[233] = 32'h00000017;
ram[234] = 32'hFFFFFF22;
ram[235] = 32'hFFFFFFE4;
ram[236] = 32'hFFFFFFE2;
ram[237] = 32'h000000FE;
ram[238] = 32'hFFFFFF4D;
ram[239] = 32'hFFFFFFD0;
ram[240] = 32'hFFFFFF6B;
ram[241] = 32'hFFFFFF8A;
ram[242] = 32'hFFFFFFCC;
ram[243] = 32'h00000010;
ram[244] = 32'hFFFFFF6D;
ram[245] = 32'hFFFFFFBE;
ram[246] = 32'h00000029;
ram[247] = 32'hFFFFFF47;
ram[248] = 32'hFFFFFFCA;
ram[249] = 32'hFFFFFF42;
ram[250] = 32'hFFFFFF8C;
ram[251] = 32'hFFFFFF25;
ram[252] = 32'h00000020;
ram[253] = 32'hFFFFFF5A;
ram[254] = 32'h00000073;
ram[255] = 32'hFFFFFF16;
ram[256] = 32'h000000D5;
ram[257] = 32'hFFFFFFF0;
ram[258] = 32'hFFFFFF3F;
ram[259] = 32'h000000A0;
ram[260] = 32'hFFFFFF7A;
ram[261] = 32'h000000BA;
ram[262] = 32'h0000006E;
ram[263] = 32'hFFFFFF17;
ram[264] = 32'hFFFFFF4D;
ram[265] = 32'hFFFFFFE3;
ram[266] = 32'hFFFFFF6C;
ram[267] = 32'hFFFFFF66;
ram[268] = 32'h000000E5;
ram[269] = 32'h0000006E;
ram[270] = 32'h000000F4;
ram[271] = 32'hFFFFFFBE;
ram[272] = 32'h000000B9;
ram[273] = 32'hFFFFFF8D;
ram[274] = 32'hFFFFFF49;
ram[275] = 32'h00000043;
ram[276] = 32'h000000ED;
ram[277] = 32'h0000005B;
ram[278] = 32'h0000008F;
ram[279] = 32'hFFFFFFBC;
ram[280] = 32'h00000048;
ram[281] = 32'hFFFFFF0E;
ram[282] = 32'h00000033;
ram[283] = 32'hFFFFFFD3;
ram[284] = 32'hFFFFFF0E;
ram[285] = 32'hFFFFFF3C;
ram[286] = 32'hFFFFFF30;
ram[287] = 32'hFFFFFFC6;
ram[288] = 32'hFFFFFF84;
ram[289] = 32'h00000014;
ram[290] = 32'hFFFFFF4A;
ram[291] = 32'hFFFFFFE0;
ram[292] = 32'h00000039;
ram[293] = 32'hFFFFFF7F;
ram[294] = 32'h00000000;
ram[295] = 32'h00000036;
ram[296] = 32'hFFFFFF98;
ram[297] = 32'hFFFFFFDC;
ram[298] = 32'h000000CE;
ram[299] = 32'h0000002D;
ram[300] = 32'hFFFFFFCB;
ram[301] = 32'hFFFFFFAC;
ram[302] = 32'hFFFFFF4A;
ram[303] = 32'h0000000C;
ram[304] = 32'h000000FB;
ram[305] = 32'h00000055;
ram[306] = 32'hFFFFFF07;
ram[307] = 32'h0000006C;
ram[308] = 32'h0000006A;
ram[309] = 32'hFFFFFF2A;
ram[310] = 32'h00000012;
ram[311] = 32'h00000060;
ram[312] = 32'h0000000A;
ram[313] = 32'hFFFFFFD3;
ram[314] = 32'hFFFFFF16;
ram[315] = 32'h0000008D;
ram[316] = 32'hFFFFFFDA;
ram[317] = 32'hFFFFFFAF;
ram[318] = 32'hFFFFFF35;
ram[319] = 32'hFFFFFFBC;
ram[320] = 32'h00000087;
ram[321] = 32'h0000007D;
ram[322] = 32'h0000003A;
ram[323] = 32'hFFFFFFAA;
ram[324] = 32'h00000023;
ram[325] = 32'hFFFFFFA8;
ram[326] = 32'hFFFFFF19;
ram[327] = 32'h00000081;
ram[328] = 32'h00000065;
ram[329] = 32'hFFFFFFDA;
ram[330] = 32'hFFFFFFAB;
ram[331] = 32'hFFFFFFF8;
ram[332] = 32'h00000093;
ram[333] = 32'hFFFFFFBB;
ram[334] = 32'hFFFFFFB7;
ram[335] = 32'h000000A5;
ram[336] = 32'h00000000;
ram[337] = 32'hFFFFFF0E;
ram[338] = 32'h00000016;
ram[339] = 32'hFFFFFF1F;
ram[340] = 32'hFFFFFF26;
ram[341] = 32'hFFFFFF59;
ram[342] = 32'h00000075;
ram[343] = 32'h00000063;
ram[344] = 32'hFFFFFF66;
ram[345] = 32'hFFFFFF93;
ram[346] = 32'h000000BD;
ram[347] = 32'hFFFFFF67;
ram[348] = 32'h000000B4;
ram[349] = 32'h00000071;
ram[350] = 32'hFFFFFF75;
ram[351] = 32'h00000067;
ram[352] = 32'h0000008E;
ram[353] = 32'hFFFFFF2F;
ram[354] = 32'h0000003F;
ram[355] = 32'h00000050;
ram[356] = 32'h00000026;
ram[357] = 32'h00000023;
ram[358] = 32'hFFFFFF0B;
ram[359] = 32'h000000D2;
ram[360] = 32'h00000083;
ram[361] = 32'h000000C0;
ram[362] = 32'h00000079;
ram[363] = 32'h00000060;
ram[364] = 32'hFFFFFF4F;
ram[365] = 32'h0000003B;
ram[366] = 32'h00000036;
ram[367] = 32'h000000FE;
ram[368] = 32'hFFFFFFB0;
ram[369] = 32'hFFFFFF95;
ram[370] = 32'hFFFFFF0B;
ram[371] = 32'h000000A8;
ram[372] = 32'hFFFFFF7D;
ram[373] = 32'hFFFFFF97;
ram[374] = 32'hFFFFFF33;
ram[375] = 32'h0000009A;
ram[376] = 32'h000000BA;
ram[377] = 32'h0000003F;
ram[378] = 32'h00000080;
ram[379] = 32'h00000069;
ram[380] = 32'hFFFFFF35;
ram[381] = 32'h0000002A;
ram[382] = 32'h00000093;
ram[383] = 32'hFFFFFF54;
ram[384] = 32'h00000023;
ram[385] = 32'h00000088;
ram[386] = 32'h00000048;
ram[387] = 32'hFFFFFF0E;
ram[388] = 32'hFFFFFFFE;
ram[389] = 32'hFFFFFF71;
ram[390] = 32'h0000004E;
ram[391] = 32'hFFFFFF75;
ram[392] = 32'hFFFFFFBE;
ram[393] = 32'h000000CC;
ram[394] = 32'hFFFFFF2C;
ram[395] = 32'h00000083;
ram[396] = 32'h0000005B;
ram[397] = 32'h0000004C;
ram[398] = 32'hFFFFFF73;
ram[399] = 32'hFFFFFF45;
ram[400] = 32'hFFFFFF07;
ram[401] = 32'h0000000B;
ram[402] = 32'h000000A6;
ram[403] = 32'h0000006C;
ram[404] = 32'h0000007E;
ram[405] = 32'hFFFFFFD5;
ram[406] = 32'h0000004A;
ram[407] = 32'hFFFFFF92;
ram[408] = 32'hFFFFFF40;
ram[409] = 32'h0000003C;
ram[410] = 32'h00000046;
ram[411] = 32'hFFFFFF49;
ram[412] = 32'h00000095;
ram[413] = 32'h000000AF;
ram[414] = 32'hFFFFFFE1;
ram[415] = 32'hFFFFFF0A;
ram[416] = 32'hFFFFFFB3;
ram[417] = 32'h0000006E;
ram[418] = 32'h000000C0;
ram[419] = 32'h00000084;
ram[420] = 32'h00000014;
ram[421] = 32'hFFFFFF48;
ram[422] = 32'h000000C1;
ram[423] = 32'hFFFFFF0D;
ram[424] = 32'h000000A7;
ram[425] = 32'h00000015;
ram[426] = 32'hFFFFFFD2;
ram[427] = 32'hFFFFFF5E;
ram[428] = 32'h000000DD;
ram[429] = 32'hFFFFFFA2;
ram[430] = 32'hFFFFFF7C;
ram[431] = 32'h00000080;
ram[432] = 32'h00000060;
ram[433] = 32'h00000090;
ram[434] = 32'hFFFFFFB4;
ram[435] = 32'h000000E0;
ram[436] = 32'hFFFFFFFC;
ram[437] = 32'h00000073;
ram[438] = 32'hFFFFFF96;
ram[439] = 32'hFFFFFF52;
ram[440] = 32'h000000CA;
ram[441] = 32'h000000FA;
ram[442] = 32'hFFFFFF61;
ram[443] = 32'h000000E7;
ram[444] = 32'h00000078;
ram[445] = 32'hFFFFFFEE;
ram[446] = 32'hFFFFFFD4;
ram[447] = 32'h0000000E;
ram[448] = 32'hFFFFFF94;
ram[449] = 32'h00000034;
ram[450] = 32'h000000C0;
ram[451] = 32'h00000087;
ram[452] = 32'h0000008E;
ram[453] = 32'hFFFFFF1A;
ram[454] = 32'h00000064;
ram[455] = 32'hFFFFFFDA;
ram[456] = 32'h00000045;
ram[457] = 32'h00000039;
ram[458] = 32'hFFFFFFE3;
ram[459] = 32'h0000005C;
ram[460] = 32'hFFFFFF9D;
ram[461] = 32'hFFFFFFFE;
ram[462] = 32'hFFFFFF8F;
ram[463] = 32'hFFFFFF62;
ram[464] = 32'h00000039;
ram[465] = 32'hFFFFFF32;
ram[466] = 32'h00000032;
ram[467] = 32'h000000E5;
ram[468] = 32'h0000008E;
ram[469] = 32'hFFFFFF7D;
ram[470] = 32'hFFFFFF5F;
ram[471] = 32'h00000071;
ram[472] = 32'h00000028;
ram[473] = 32'h00000098;
ram[474] = 32'hFFFFFF4B;
ram[475] = 32'hFFFFFF06;
ram[476] = 32'h00000069;
ram[477] = 32'h00000079;
ram[478] = 32'h000000A2;
ram[479] = 32'h00000037;
ram[480] = 32'h000000C5;
ram[481] = 32'h0000009F;
ram[482] = 32'hFFFFFF57;
ram[483] = 32'hFFFFFFF0;
ram[484] = 32'h000000BA;
ram[485] = 32'h000000FD;
ram[486] = 32'h000000BA;
ram[487] = 32'h00000075;
ram[488] = 32'h0000003B;
ram[489] = 32'hFFFFFFD8;
ram[490] = 32'h000000E3;
ram[491] = 32'hFFFFFF6E;
ram[492] = 32'h0000000B;
ram[493] = 32'hFFFFFF9C;
ram[494] = 32'h00000019;
ram[495] = 32'h000000BB;
ram[496] = 32'hFFFFFF92;
ram[497] = 32'hFFFFFF39;
ram[498] = 32'h000000FE;
ram[499] = 32'h0000004D;
ram[500] = 32'h00000070;
ram[501] = 32'h0000008F;
ram[502] = 32'hFFFFFF9A;
ram[503] = 32'hFFFFFF4D;
ram[504] = 32'hFFFFFFE9;
ram[505] = 32'hFFFFFF7D;
ram[506] = 32'h00000000;
ram[507] = 32'h00000071;
ram[508] = 32'h000000D6;
ram[509] = 32'hFFFFFF05;
ram[510] = 32'hFFFFFF58;
ram[511] = 32'hFFFFFF84;

end

  //-- Lectura de la memoria
  always @ * begin
    if (rw == 1)
    data_out <= ram[addr];
  end

  //-- Escritura en la memoria



  always @ * begin
    if (rw == 0)
     ram[addr] <= data_in;
  end




endmodule
